`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.08.2023 21:02:18
// Design Name: 
// Module Name: otfs
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module otfs(        xin1, xin2, xin3, xin4, xin5, xin6, xin7, xin8, xin9, xin10, xin11, xin12, xin13, xin14, xin15, xin16, xin17, xin18, xin19, xin20, xin21, xin22, xin23, xin24, xin25, xin26, xin27, xin28, xin29, xin30, xin31, xin32, xin33, xin34, xin35, xin36, xin37, xin38, xin39, xin40, xin41, xin42, xin43, xin44, xin45, xin46, xin47, xin48, xin49, xin50, xin51, xin52, xin53, xin54, xin55, xin56, xin57, xin58, xin59, xin60, xin61, xin62, xin63, xin64, xin65, xin66, xin67, xin68, xin69, xin70, xin71, xin72, xin73, xin74, xin75, xin76, xin77, xin78, xin79, xin80, xin81, xin82, xin83, xin84, xin85, xin86, xin87, xin88, xin89, xin90, xin91, xin92, xin93, xin94, xin95, xin96, xin97, xin98, xin99, xin100, xin101, xin102, xin103, xin104, xin105, xin106, xin107, xin108, xin109, xin110, xin111, xin112, xin113, xin114, xin115, xin116, xin117, xin118, xin119, xin120, xin121, xin122, xin123, xin124, xin125, xin126, xin127, xin128, xin129, xin130, xin131, xin132, xin133, xin134, xin135, xin136, xin137, xin138, xin139, xin140, xin141, xin142, xin143, xin144, xin145, xin146, xin147, xin148, xin149, xin150, xin151, xin152, xin153, xin154, xin155, xin156, xin157, xin158, xin159, xin160, xin161, xin162, xin163, xin164, xin165, xin166, xin167, xin168, xin169, xin170, xin171, xin172, xin173, xin174, xin175, xin176, xin177, xin178, xin179, xin180, xin181, xin182, xin183, xin184, xin185, xin186, xin187, xin188, xin189, xin190, xin191, xin192, xin193, xin194, xin195, xin196, xin197, xin198, xin199, xin200, xin201, xin202, xin203, xin204, xin205, xin206, xin207, xin208, xin209, xin210, xin211, xin212, xin213, xin214, xin215, xin216, xin217, xin218, xin219, xin220, xin221, xin222, xin223, xin224, xin225, xin226, xin227, xin228, xin229, xin230, xin231, xin232, xin233, xin234, xin235, xin236, xin237, xin238, xin239, xin240, xin241, xin242, xin243, xin244, xin245, xin246, xin247, xin248, xin249, xin250, xin251, xin252, xin253, xin254, xin255, xin256,
                    yin1, yin2, yin3, yin4, yin5, yin6, yin7, yin8, yin9, yin10, yin11, yin12, yin13, yin14, yin15, yin16, yin17, yin18, yin19, yin20, yin21, yin22, yin23, yin24, yin25, yin26, yin27, yin28, yin29, yin30, yin31, yin32, yin33, yin34, yin35, yin36, yin37, yin38, yin39, yin40, yin41, yin42, yin43, yin44, yin45, yin46, yin47, yin48, yin49, yin50, yin51, yin52, yin53, yin54, yin55, yin56, yin57, yin58, yin59, yin60, yin61, yin62, yin63, yin64, yin65, yin66, yin67, yin68, yin69, yin70, yin71, yin72, yin73, yin74, yin75, yin76, yin77, yin78, yin79, yin80, yin81, yin82, yin83, yin84, yin85, yin86, yin87, yin88, yin89, yin90, yin91, yin92, yin93, yin94, yin95, yin96, yin97, yin98, yin99, yin100, yin101, yin102, yin103, yin104, yin105, yin106, yin107, yin108, yin109, yin110, yin111, yin112, yin113, yin114, yin115, yin116, yin117, yin118, yin119, yin120, yin121, yin122, yin123, yin124, yin125, yin126, yin127, yin128, yin129, yin130, yin131, yin132, yin133, yin134, yin135, yin136, yin137, yin138, yin139, yin140, yin141, yin142, yin143, yin144, yin145, yin146, yin147, yin148, yin149, yin150, yin151, yin152, yin153, yin154, yin155, yin156, yin157, yin158, yin159, yin160, yin161, yin162, yin163, yin164, yin165, yin166, yin167, yin168, yin169, yin170, yin171, yin172, yin173, yin174, yin175, yin176, yin177, yin178, yin179, yin180, yin181, yin182, yin183, yin184, yin185, yin186, yin187, yin188, yin189, yin190, yin191, yin192, yin193, yin194, yin195, yin196, yin197, yin198, yin199, yin200, yin201, yin202, yin203, yin204, yin205, yin206, yin207, yin208, yin209, yin210, yin211, yin212, yin213, yin214, yin215, yin216, yin217, yin218, yin219, yin220, yin221, yin222, yin223, yin224, yin225, yin226, yin227, yin228, yin229, yin230, yin231, yin232, yin233, yin234, yin235, yin236, yin237, yin238, yin239, yin240, yin241, yin242, yin243, yin244, yin245, yin246, yin247, yin248, yin249, yin250, yin251, yin252, yin253, yin254, yin255, yin256,
                    clock,
                    xout1, xout2, xout3, xout4, xout5, xout6, xout7, xout8, xout9, xout10, xout11, xout12, xout13, xout14, xout15, xout16, xout17, xout18, xout19, xout20, xout21, xout22, xout23, xout24, xout25, xout26, xout27, xout28, xout29, xout30, xout31, xout32, xout33, xout34, xout35, xout36, xout37, xout38, xout39, xout40, xout41, xout42, xout43, xout44, xout45, xout46, xout47, xout48, xout49, xout50, xout51, xout52, xout53, xout54, xout55, xout56, xout57, xout58, xout59, xout60, xout61, xout62, xout63, xout64, xout65, xout66, xout67, xout68, xout69, xout70, xout71, xout72, xout73, xout74, xout75, xout76, xout77, xout78, xout79, xout80, xout81, xout82, xout83, xout84, xout85, xout86, xout87, xout88, xout89, xout90, xout91, xout92, xout93, xout94, xout95, xout96, xout97, xout98, xout99, xout100, xout101, xout102, xout103, xout104, xout105, xout106, xout107, xout108, xout109, xout110, xout111, xout112, xout113, xout114, xout115, xout116, xout117, xout118, xout119, xout120, xout121, xout122, xout123, xout124, xout125, xout126, xout127, xout128, xout129, xout130, xout131, xout132, xout133, xout134, xout135, xout136, xout137, xout138, xout139, xout140, xout141, xout142, xout143, xout144, xout145, xout146, xout147, xout148, xout149, xout150, xout151, xout152, xout153, xout154, xout155, xout156, xout157, xout158, xout159, xout160, xout161, xout162, xout163, xout164, xout165, xout166, xout167, xout168, xout169, xout170, xout171, xout172, xout173, xout174, xout175, xout176, xout177, xout178, xout179, xout180, xout181, xout182, xout183, xout184, xout185, xout186, xout187, xout188, xout189, xout190, xout191, xout192, xout193, xout194, xout195, xout196, xout197, xout198, xout199, xout200, xout201, xout202, xout203, xout204, xout205, xout206, xout207, xout208, xout209, xout210, xout211, xout212, xout213, xout214, xout215, xout216, xout217, xout218, xout219, xout220, xout221, xout222, xout223, xout224, xout225, xout226, xout227, xout228, xout229, xout230, xout231, xout232, xout233, xout234, xout235, xout236, xout237, xout238, xout239, xout240, xout241, xout242, xout243, xout244, xout245, xout246, xout247, xout248, xout249, xout250, xout251, xout252, xout253, xout254, xout255, xout256,
                    yout1, yout2, yout3, yout4, yout5, yout6, yout7, yout8, yout9, yout10, yout11, yout12, yout13, yout14, yout15, yout16, yout17, yout18, yout19, yout20, yout21, yout22, yout23, yout24, yout25, yout26, yout27, yout28, yout29, yout30, yout31, yout32, yout33, yout34, yout35, yout36, yout37, yout38, yout39, yout40, yout41, yout42, yout43, yout44, yout45, yout46, yout47, yout48, yout49, yout50, yout51, yout52, yout53, yout54, yout55, yout56, yout57, yout58, yout59, yout60, yout61, yout62, yout63, yout64, yout65, yout66, yout67, yout68, yout69, yout70, yout71, yout72, yout73, yout74, yout75, yout76, yout77, yout78, yout79, yout80, yout81, yout82, yout83, yout84, yout85, yout86, yout87, yout88, yout89, yout90, yout91, yout92, yout93, yout94, yout95, yout96, yout97, yout98, yout99, yout100, yout101, yout102, yout103, yout104, yout105, yout106, yout107, yout108, yout109, yout110, yout111, yout112, yout113, yout114, yout115, yout116, yout117, yout118, yout119, yout120, yout121, yout122, yout123, yout124, yout125, yout126, yout127, yout128, yout129, yout130, yout131, yout132, yout133, yout134, yout135, yout136, yout137, yout138, yout139, yout140, yout141, yout142, yout143, yout144, yout145, yout146, yout147, yout148, yout149, yout150, yout151, yout152, yout153, yout154, yout155, yout156, yout157, yout158, yout159, yout160, yout161, yout162, yout163, yout164, yout165, yout166, yout167, yout168, yout169, yout170, yout171, yout172, yout173, yout174, yout175, yout176, yout177, yout178, yout179, yout180, yout181, yout182, yout183, yout184, yout185, yout186, yout187, yout188, yout189, yout190, yout191, yout192, yout193, yout194, yout195, yout196, yout197, yout198, yout199, yout200, yout201, yout202, yout203, yout204, yout205, yout206, yout207, yout208, yout209, yout210, yout211, yout212, yout213, yout214, yout215, yout216, yout217, yout218, yout219, yout220, yout221, yout222, yout223, yout224, yout225, yout226, yout227, yout228, yout229, yout230, yout231, yout232, yout233, yout234, yout235, yout236, yout237, yout238, yout239, yout240, yout241, yout242, yout243, yout244, yout245, yout246, yout247, yout248, yout249, yout250, yout251, yout252, yout253, yout254, yout255, yout256
            );

    
input signed [15:0] xin1;
input signed [15:0] xin2;
input signed [15:0] xin3;
input signed [15:0] xin4;
input signed [15:0] xin5;
input signed [15:0] xin6;
input signed [15:0] xin7;
input signed [15:0] xin8;
input signed [15:0] xin9;
input signed [15:0] xin10;
input signed [15:0] xin11;
input signed [15:0] xin12;
input signed [15:0] xin13;
input signed [15:0] xin14;
input signed [15:0] xin15;
input signed [15:0] xin16;
input signed [15:0] xin17;
input signed [15:0] xin18;
input signed [15:0] xin19;
input signed [15:0] xin20;
input signed [15:0] xin21;
input signed [15:0] xin22;
input signed [15:0] xin23;
input signed [15:0] xin24;
input signed [15:0] xin25;
input signed [15:0] xin26;
input signed [15:0] xin27;
input signed [15:0] xin28;
input signed [15:0] xin29;
input signed [15:0] xin30;
input signed [15:0] xin31;
input signed [15:0] xin32;
input signed [15:0] xin33;
input signed [15:0] xin34;
input signed [15:0] xin35;
input signed [15:0] xin36;
input signed [15:0] xin37;
input signed [15:0] xin38;
input signed [15:0] xin39;
input signed [15:0] xin40;
input signed [15:0] xin41;
input signed [15:0] xin42;
input signed [15:0] xin43;
input signed [15:0] xin44;
input signed [15:0] xin45;
input signed [15:0] xin46;
input signed [15:0] xin47;
input signed [15:0] xin48;
input signed [15:0] xin49;
input signed [15:0] xin50;
input signed [15:0] xin51;
input signed [15:0] xin52;
input signed [15:0] xin53;
input signed [15:0] xin54;
input signed [15:0] xin55;
input signed [15:0] xin56;
input signed [15:0] xin57;
input signed [15:0] xin58;
input signed [15:0] xin59;
input signed [15:0] xin60;
input signed [15:0] xin61;
input signed [15:0] xin62;
input signed [15:0] xin63;
input signed [15:0] xin64;
input signed [15:0] xin65;
input signed [15:0] xin66;
input signed [15:0] xin67;
input signed [15:0] xin68;
input signed [15:0] xin69;
input signed [15:0] xin70;
input signed [15:0] xin71;
input signed [15:0] xin72;
input signed [15:0] xin73;
input signed [15:0] xin74;
input signed [15:0] xin75;
input signed [15:0] xin76;
input signed [15:0] xin77;
input signed [15:0] xin78;
input signed [15:0] xin79;
input signed [15:0] xin80;
input signed [15:0] xin81;
input signed [15:0] xin82;
input signed [15:0] xin83;
input signed [15:0] xin84;
input signed [15:0] xin85;
input signed [15:0] xin86;
input signed [15:0] xin87;
input signed [15:0] xin88;
input signed [15:0] xin89;
input signed [15:0] xin90;
input signed [15:0] xin91;
input signed [15:0] xin92;
input signed [15:0] xin93;
input signed [15:0] xin94;
input signed [15:0] xin95;
input signed [15:0] xin96;
input signed [15:0] xin97;
input signed [15:0] xin98;
input signed [15:0] xin99;
input signed [15:0] xin100;
input signed [15:0] xin101;
input signed [15:0] xin102;
input signed [15:0] xin103;
input signed [15:0] xin104;
input signed [15:0] xin105;
input signed [15:0] xin106;
input signed [15:0] xin107;
input signed [15:0] xin108;
input signed [15:0] xin109;
input signed [15:0] xin110;
input signed [15:0] xin111;
input signed [15:0] xin112;
input signed [15:0] xin113;
input signed [15:0] xin114;
input signed [15:0] xin115;
input signed [15:0] xin116;
input signed [15:0] xin117;
input signed [15:0] xin118;
input signed [15:0] xin119;
input signed [15:0] xin120;
input signed [15:0] xin121;
input signed [15:0] xin122;
input signed [15:0] xin123;
input signed [15:0] xin124;
input signed [15:0] xin125;
input signed [15:0] xin126;
input signed [15:0] xin127;
input signed [15:0] xin128;
input signed [15:0] xin129;
input signed [15:0] xin130;
input signed [15:0] xin131;
input signed [15:0] xin132;
input signed [15:0] xin133;
input signed [15:0] xin134;
input signed [15:0] xin135;
input signed [15:0] xin136;
input signed [15:0] xin137;
input signed [15:0] xin138;
input signed [15:0] xin139;
input signed [15:0] xin140;
input signed [15:0] xin141;
input signed [15:0] xin142;
input signed [15:0] xin143;
input signed [15:0] xin144;
input signed [15:0] xin145;
input signed [15:0] xin146;
input signed [15:0] xin147;
input signed [15:0] xin148;
input signed [15:0] xin149;
input signed [15:0] xin150;
input signed [15:0] xin151;
input signed [15:0] xin152;
input signed [15:0] xin153;
input signed [15:0] xin154;
input signed [15:0] xin155;
input signed [15:0] xin156;
input signed [15:0] xin157;
input signed [15:0] xin158;
input signed [15:0] xin159;
input signed [15:0] xin160;
input signed [15:0] xin161;
input signed [15:0] xin162;
input signed [15:0] xin163;
input signed [15:0] xin164;
input signed [15:0] xin165;
input signed [15:0] xin166;
input signed [15:0] xin167;
input signed [15:0] xin168;
input signed [15:0] xin169;
input signed [15:0] xin170;
input signed [15:0] xin171;
input signed [15:0] xin172;
input signed [15:0] xin173;
input signed [15:0] xin174;
input signed [15:0] xin175;
input signed [15:0] xin176;
input signed [15:0] xin177;
input signed [15:0] xin178;
input signed [15:0] xin179;
input signed [15:0] xin180;
input signed [15:0] xin181;
input signed [15:0] xin182;
input signed [15:0] xin183;
input signed [15:0] xin184;
input signed [15:0] xin185;
input signed [15:0] xin186;
input signed [15:0] xin187;
input signed [15:0] xin188;
input signed [15:0] xin189;
input signed [15:0] xin190;
input signed [15:0] xin191;
input signed [15:0] xin192;
input signed [15:0] xin193;
input signed [15:0] xin194;
input signed [15:0] xin195;
input signed [15:0] xin196;
input signed [15:0] xin197;
input signed [15:0] xin198;
input signed [15:0] xin199;
input signed [15:0] xin200;
input signed [15:0] xin201;
input signed [15:0] xin202;
input signed [15:0] xin203;
input signed [15:0] xin204;
input signed [15:0] xin205;
input signed [15:0] xin206;
input signed [15:0] xin207;
input signed [15:0] xin208;
input signed [15:0] xin209;
input signed [15:0] xin210;
input signed [15:0] xin211;
input signed [15:0] xin212;
input signed [15:0] xin213;
input signed [15:0] xin214;
input signed [15:0] xin215;
input signed [15:0] xin216;
input signed [15:0] xin217;
input signed [15:0] xin218;
input signed [15:0] xin219;
input signed [15:0] xin220;
input signed [15:0] xin221;
input signed [15:0] xin222;
input signed [15:0] xin223;
input signed [15:0] xin224;
input signed [15:0] xin225;
input signed [15:0] xin226;
input signed [15:0] xin227;
input signed [15:0] xin228;
input signed [15:0] xin229;
input signed [15:0] xin230;
input signed [15:0] xin231;
input signed [15:0] xin232;
input signed [15:0] xin233;
input signed [15:0] xin234;
input signed [15:0] xin235;
input signed [15:0] xin236;
input signed [15:0] xin237;
input signed [15:0] xin238;
input signed [15:0] xin239;
input signed [15:0] xin240;
input signed [15:0] xin241;
input signed [15:0] xin242;
input signed [15:0] xin243;
input signed [15:0] xin244;
input signed [15:0] xin245;
input signed [15:0] xin246;
input signed [15:0] xin247;
input signed [15:0] xin248;
input signed [15:0] xin249;
input signed [15:0] xin250;
input signed [15:0] xin251;
input signed [15:0] xin252;
input signed [15:0] xin253;
input signed [15:0] xin254;
input signed [15:0] xin255;
input signed [15:0] xin256;

input signed [15:0] yin1;
input signed [15:0] yin2;
input signed [15:0] yin3;
input signed [15:0] yin4;
input signed [15:0] yin5;
input signed [15:0] yin6;
input signed [15:0] yin7;
input signed [15:0] yin8;
input signed [15:0] yin9;
input signed [15:0] yin10;
input signed [15:0] yin11;
input signed [15:0] yin12;
input signed [15:0] yin13;
input signed [15:0] yin14;
input signed [15:0] yin15;
input signed [15:0] yin16;
input signed [15:0] yin17;
input signed [15:0] yin18;
input signed [15:0] yin19;
input signed [15:0] yin20;
input signed [15:0] yin21;
input signed [15:0] yin22;
input signed [15:0] yin23;
input signed [15:0] yin24;
input signed [15:0] yin25;
input signed [15:0] yin26;
input signed [15:0] yin27;
input signed [15:0] yin28;
input signed [15:0] yin29;
input signed [15:0] yin30;
input signed [15:0] yin31;
input signed [15:0] yin32;
input signed [15:0] yin33;
input signed [15:0] yin34;
input signed [15:0] yin35;
input signed [15:0] yin36;
input signed [15:0] yin37;
input signed [15:0] yin38;
input signed [15:0] yin39;
input signed [15:0] yin40;
input signed [15:0] yin41;
input signed [15:0] yin42;
input signed [15:0] yin43;
input signed [15:0] yin44;
input signed [15:0] yin45;
input signed [15:0] yin46;
input signed [15:0] yin47;
input signed [15:0] yin48;
input signed [15:0] yin49;
input signed [15:0] yin50;
input signed [15:0] yin51;
input signed [15:0] yin52;
input signed [15:0] yin53;
input signed [15:0] yin54;
input signed [15:0] yin55;
input signed [15:0] yin56;
input signed [15:0] yin57;
input signed [15:0] yin58;
input signed [15:0] yin59;
input signed [15:0] yin60;
input signed [15:0] yin61;
input signed [15:0] yin62;
input signed [15:0] yin63;
input signed [15:0] yin64;
input signed [15:0] yin65;
input signed [15:0] yin66;
input signed [15:0] yin67;
input signed [15:0] yin68;
input signed [15:0] yin69;
input signed [15:0] yin70;
input signed [15:0] yin71;
input signed [15:0] yin72;
input signed [15:0] yin73;
input signed [15:0] yin74;
input signed [15:0] yin75;
input signed [15:0] yin76;
input signed [15:0] yin77;
input signed [15:0] yin78;
input signed [15:0] yin79;
input signed [15:0] yin80;
input signed [15:0] yin81;
input signed [15:0] yin82;
input signed [15:0] yin83;
input signed [15:0] yin84;
input signed [15:0] yin85;
input signed [15:0] yin86;
input signed [15:0] yin87;
input signed [15:0] yin88;
input signed [15:0] yin89;
input signed [15:0] yin90;
input signed [15:0] yin91;
input signed [15:0] yin92;
input signed [15:0] yin93;
input signed [15:0] yin94;
input signed [15:0] yin95;
input signed [15:0] yin96;
input signed [15:0] yin97;
input signed [15:0] yin98;
input signed [15:0] yin99;
input signed [15:0] yin100;
input signed [15:0] yin101;
input signed [15:0] yin102;
input signed [15:0] yin103;
input signed [15:0] yin104;
input signed [15:0] yin105;
input signed [15:0] yin106;
input signed [15:0] yin107;
input signed [15:0] yin108;
input signed [15:0] yin109;
input signed [15:0] yin110;
input signed [15:0] yin111;
input signed [15:0] yin112;
input signed [15:0] yin113;
input signed [15:0] yin114;
input signed [15:0] yin115;
input signed [15:0] yin116;
input signed [15:0] yin117;
input signed [15:0] yin118;
input signed [15:0] yin119;
input signed [15:0] yin120;
input signed [15:0] yin121;
input signed [15:0] yin122;
input signed [15:0] yin123;
input signed [15:0] yin124;
input signed [15:0] yin125;
input signed [15:0] yin126;
input signed [15:0] yin127;
input signed [15:0] yin128;
input signed [15:0] yin129;
input signed [15:0] yin130;
input signed [15:0] yin131;
input signed [15:0] yin132;
input signed [15:0] yin133;
input signed [15:0] yin134;
input signed [15:0] yin135;
input signed [15:0] yin136;
input signed [15:0] yin137;
input signed [15:0] yin138;
input signed [15:0] yin139;
input signed [15:0] yin140;
input signed [15:0] yin141;
input signed [15:0] yin142;
input signed [15:0] yin143;
input signed [15:0] yin144;
input signed [15:0] yin145;
input signed [15:0] yin146;
input signed [15:0] yin147;
input signed [15:0] yin148;
input signed [15:0] yin149;
input signed [15:0] yin150;
input signed [15:0] yin151;
input signed [15:0] yin152;
input signed [15:0] yin153;
input signed [15:0] yin154;
input signed [15:0] yin155;
input signed [15:0] yin156;
input signed [15:0] yin157;
input signed [15:0] yin158;
input signed [15:0] yin159;
input signed [15:0] yin160;
input signed [15:0] yin161;
input signed [15:0] yin162;
input signed [15:0] yin163;
input signed [15:0] yin164;
input signed [15:0] yin165;
input signed [15:0] yin166;
input signed [15:0] yin167;
input signed [15:0] yin168;
input signed [15:0] yin169;
input signed [15:0] yin170;
input signed [15:0] yin171;
input signed [15:0] yin172;
input signed [15:0] yin173;
input signed [15:0] yin174;
input signed [15:0] yin175;
input signed [15:0] yin176;
input signed [15:0] yin177;
input signed [15:0] yin178;
input signed [15:0] yin179;
input signed [15:0] yin180;
input signed [15:0] yin181;
input signed [15:0] yin182;
input signed [15:0] yin183;
input signed [15:0] yin184;
input signed [15:0] yin185;
input signed [15:0] yin186;
input signed [15:0] yin187;
input signed [15:0] yin188;
input signed [15:0] yin189;
input signed [15:0] yin190;
input signed [15:0] yin191;
input signed [15:0] yin192;
input signed [15:0] yin193;
input signed [15:0] yin194;
input signed [15:0] yin195;
input signed [15:0] yin196;
input signed [15:0] yin197;
input signed [15:0] yin198;
input signed [15:0] yin199;
input signed [15:0] yin200;
input signed [15:0] yin201;
input signed [15:0] yin202;
input signed [15:0] yin203;
input signed [15:0] yin204;
input signed [15:0] yin205;
input signed [15:0] yin206;
input signed [15:0] yin207;
input signed [15:0] yin208;
input signed [15:0] yin209;
input signed [15:0] yin210;
input signed [15:0] yin211;
input signed [15:0] yin212;
input signed [15:0] yin213;
input signed [15:0] yin214;
input signed [15:0] yin215;
input signed [15:0] yin216;
input signed [15:0] yin217;
input signed [15:0] yin218;
input signed [15:0] yin219;
input signed [15:0] yin220;
input signed [15:0] yin221;
input signed [15:0] yin222;
input signed [15:0] yin223;
input signed [15:0] yin224;
input signed [15:0] yin225;
input signed [15:0] yin226;
input signed [15:0] yin227;
input signed [15:0] yin228;
input signed [15:0] yin229;
input signed [15:0] yin230;
input signed [15:0] yin231;
input signed [15:0] yin232;
input signed [15:0] yin233;
input signed [15:0] yin234;
input signed [15:0] yin235;
input signed [15:0] yin236;
input signed [15:0] yin237;
input signed [15:0] yin238;
input signed [15:0] yin239;
input signed [15:0] yin240;
input signed [15:0] yin241;
input signed [15:0] yin242;
input signed [15:0] yin243;
input signed [15:0] yin244;
input signed [15:0] yin245;
input signed [15:0] yin246;
input signed [15:0] yin247;
input signed [15:0] yin248;
input signed [15:0] yin249;
input signed [15:0] yin250;
input signed [15:0] yin251;
input signed [15:0] yin252;
input signed [15:0] yin253;
input signed [15:0] yin254;
input signed [15:0] yin255;
input signed [15:0] yin256;

input clock;

output signed [15:0] xout1;
output signed [15:0] xout2;
output signed [15:0] xout3;
output signed [15:0] xout4;
output signed [15:0] xout5;
output signed [15:0] xout6;
output signed [15:0] xout7;
output signed [15:0] xout8;
output signed [15:0] xout9;
output signed [15:0] xout10;
output signed [15:0] xout11;
output signed [15:0] xout12;
output signed [15:0] xout13;
output signed [15:0] xout14;
output signed [15:0] xout15;
output signed [15:0] xout16;
output signed [15:0] xout17;
output signed [15:0] xout18;
output signed [15:0] xout19;
output signed [15:0] xout20;
output signed [15:0] xout21;
output signed [15:0] xout22;
output signed [15:0] xout23;
output signed [15:0] xout24;
output signed [15:0] xout25;
output signed [15:0] xout26;
output signed [15:0] xout27;
output signed [15:0] xout28;
output signed [15:0] xout29;
output signed [15:0] xout30;
output signed [15:0] xout31;
output signed [15:0] xout32;
output signed [15:0] xout33;
output signed [15:0] xout34;
output signed [15:0] xout35;
output signed [15:0] xout36;
output signed [15:0] xout37;
output signed [15:0] xout38;
output signed [15:0] xout39;
output signed [15:0] xout40;
output signed [15:0] xout41;
output signed [15:0] xout42;
output signed [15:0] xout43;
output signed [15:0] xout44;
output signed [15:0] xout45;
output signed [15:0] xout46;
output signed [15:0] xout47;
output signed [15:0] xout48;
output signed [15:0] xout49;
output signed [15:0] xout50;
output signed [15:0] xout51;
output signed [15:0] xout52;
output signed [15:0] xout53;
output signed [15:0] xout54;
output signed [15:0] xout55;
output signed [15:0] xout56;
output signed [15:0] xout57;
output signed [15:0] xout58;
output signed [15:0] xout59;
output signed [15:0] xout60;
output signed [15:0] xout61;
output signed [15:0] xout62;
output signed [15:0] xout63;
output signed [15:0] xout64;
output signed [15:0] xout65;
output signed [15:0] xout66;
output signed [15:0] xout67;
output signed [15:0] xout68;
output signed [15:0] xout69;
output signed [15:0] xout70;
output signed [15:0] xout71;
output signed [15:0] xout72;
output signed [15:0] xout73;
output signed [15:0] xout74;
output signed [15:0] xout75;
output signed [15:0] xout76;
output signed [15:0] xout77;
output signed [15:0] xout78;
output signed [15:0] xout79;
output signed [15:0] xout80;
output signed [15:0] xout81;
output signed [15:0] xout82;
output signed [15:0] xout83;
output signed [15:0] xout84;
output signed [15:0] xout85;
output signed [15:0] xout86;
output signed [15:0] xout87;
output signed [15:0] xout88;
output signed [15:0] xout89;
output signed [15:0] xout90;
output signed [15:0] xout91;
output signed [15:0] xout92;
output signed [15:0] xout93;
output signed [15:0] xout94;
output signed [15:0] xout95;
output signed [15:0] xout96;
output signed [15:0] xout97;
output signed [15:0] xout98;
output signed [15:0] xout99;
output signed [15:0] xout100;
output signed [15:0] xout101;
output signed [15:0] xout102;
output signed [15:0] xout103;
output signed [15:0] xout104;
output signed [15:0] xout105;
output signed [15:0] xout106;
output signed [15:0] xout107;
output signed [15:0] xout108;
output signed [15:0] xout109;
output signed [15:0] xout110;
output signed [15:0] xout111;
output signed [15:0] xout112;
output signed [15:0] xout113;
output signed [15:0] xout114;
output signed [15:0] xout115;
output signed [15:0] xout116;
output signed [15:0] xout117;
output signed [15:0] xout118;
output signed [15:0] xout119;
output signed [15:0] xout120;
output signed [15:0] xout121;
output signed [15:0] xout122;
output signed [15:0] xout123;
output signed [15:0] xout124;
output signed [15:0] xout125;
output signed [15:0] xout126;
output signed [15:0] xout127;
output signed [15:0] xout128;
output signed [15:0] xout129;
output signed [15:0] xout130;
output signed [15:0] xout131;
output signed [15:0] xout132;
output signed [15:0] xout133;
output signed [15:0] xout134;
output signed [15:0] xout135;
output signed [15:0] xout136;
output signed [15:0] xout137;
output signed [15:0] xout138;
output signed [15:0] xout139;
output signed [15:0] xout140;
output signed [15:0] xout141;
output signed [15:0] xout142;
output signed [15:0] xout143;
output signed [15:0] xout144;
output signed [15:0] xout145;
output signed [15:0] xout146;
output signed [15:0] xout147;
output signed [15:0] xout148;
output signed [15:0] xout149;
output signed [15:0] xout150;
output signed [15:0] xout151;
output signed [15:0] xout152;
output signed [15:0] xout153;
output signed [15:0] xout154;
output signed [15:0] xout155;
output signed [15:0] xout156;
output signed [15:0] xout157;
output signed [15:0] xout158;
output signed [15:0] xout159;
output signed [15:0] xout160;
output signed [15:0] xout161;
output signed [15:0] xout162;
output signed [15:0] xout163;
output signed [15:0] xout164;
output signed [15:0] xout165;
output signed [15:0] xout166;
output signed [15:0] xout167;
output signed [15:0] xout168;
output signed [15:0] xout169;
output signed [15:0] xout170;
output signed [15:0] xout171;
output signed [15:0] xout172;
output signed [15:0] xout173;
output signed [15:0] xout174;
output signed [15:0] xout175;
output signed [15:0] xout176;
output signed [15:0] xout177;
output signed [15:0] xout178;
output signed [15:0] xout179;
output signed [15:0] xout180;
output signed [15:0] xout181;
output signed [15:0] xout182;
output signed [15:0] xout183;
output signed [15:0] xout184;
output signed [15:0] xout185;
output signed [15:0] xout186;
output signed [15:0] xout187;
output signed [15:0] xout188;
output signed [15:0] xout189;
output signed [15:0] xout190;
output signed [15:0] xout191;
output signed [15:0] xout192;
output signed [15:0] xout193;
output signed [15:0] xout194;
output signed [15:0] xout195;
output signed [15:0] xout196;
output signed [15:0] xout197;
output signed [15:0] xout198;
output signed [15:0] xout199;
output signed [15:0] xout200;
output signed [15:0] xout201;
output signed [15:0] xout202;
output signed [15:0] xout203;
output signed [15:0] xout204;
output signed [15:0] xout205;
output signed [15:0] xout206;
output signed [15:0] xout207;
output signed [15:0] xout208;
output signed [15:0] xout209;
output signed [15:0] xout210;
output signed [15:0] xout211;
output signed [15:0] xout212;
output signed [15:0] xout213;
output signed [15:0] xout214;
output signed [15:0] xout215;
output signed [15:0] xout216;
output signed [15:0] xout217;
output signed [15:0] xout218;
output signed [15:0] xout219;
output signed [15:0] xout220;
output signed [15:0] xout221;
output signed [15:0] xout222;
output signed [15:0] xout223;
output signed [15:0] xout224;
output signed [15:0] xout225;
output signed [15:0] xout226;
output signed [15:0] xout227;
output signed [15:0] xout228;
output signed [15:0] xout229;
output signed [15:0] xout230;
output signed [15:0] xout231;
output signed [15:0] xout232;
output signed [15:0] xout233;
output signed [15:0] xout234;
output signed [15:0] xout235;
output signed [15:0] xout236;
output signed [15:0] xout237;
output signed [15:0] xout238;
output signed [15:0] xout239;
output signed [15:0] xout240;
output signed [15:0] xout241;
output signed [15:0] xout242;
output signed [15:0] xout243;
output signed [15:0] xout244;
output signed [15:0] xout245;
output signed [15:0] xout246;
output signed [15:0] xout247;
output signed [15:0] xout248;
output signed [15:0] xout249;
output signed [15:0] xout250;
output signed [15:0] xout251;
output signed [15:0] xout252;
output signed [15:0] xout253;
output signed [15:0] xout254;
output signed [15:0] xout255;
output signed [15:0] xout256;

output signed [15:0] yout1;
output signed [15:0] yout2;
output signed [15:0] yout3;
output signed [15:0] yout4;
output signed [15:0] yout5;
output signed [15:0] yout6;
output signed [15:0] yout7;
output signed [15:0] yout8;
output signed [15:0] yout9;
output signed [15:0] yout10;
output signed [15:0] yout11;
output signed [15:0] yout12;
output signed [15:0] yout13;
output signed [15:0] yout14;
output signed [15:0] yout15;
output signed [15:0] yout16;
output signed [15:0] yout17;
output signed [15:0] yout18;
output signed [15:0] yout19;
output signed [15:0] yout20;
output signed [15:0] yout21;
output signed [15:0] yout22;
output signed [15:0] yout23;
output signed [15:0] yout24;
output signed [15:0] yout25;
output signed [15:0] yout26;
output signed [15:0] yout27;
output signed [15:0] yout28;
output signed [15:0] yout29;
output signed [15:0] yout30;
output signed [15:0] yout31;
output signed [15:0] yout32;
output signed [15:0] yout33;
output signed [15:0] yout34;
output signed [15:0] yout35;
output signed [15:0] yout36;
output signed [15:0] yout37;
output signed [15:0] yout38;
output signed [15:0] yout39;
output signed [15:0] yout40;
output signed [15:0] yout41;
output signed [15:0] yout42;
output signed [15:0] yout43;
output signed [15:0] yout44;
output signed [15:0] yout45;
output signed [15:0] yout46;
output signed [15:0] yout47;
output signed [15:0] yout48;
output signed [15:0] yout49;
output signed [15:0] yout50;
output signed [15:0] yout51;
output signed [15:0] yout52;
output signed [15:0] yout53;
output signed [15:0] yout54;
output signed [15:0] yout55;
output signed [15:0] yout56;
output signed [15:0] yout57;
output signed [15:0] yout58;
output signed [15:0] yout59;
output signed [15:0] yout60;
output signed [15:0] yout61;
output signed [15:0] yout62;
output signed [15:0] yout63;
output signed [15:0] yout64;
output signed [15:0] yout65;
output signed [15:0] yout66;
output signed [15:0] yout67;
output signed [15:0] yout68;
output signed [15:0] yout69;
output signed [15:0] yout70;
output signed [15:0] yout71;
output signed [15:0] yout72;
output signed [15:0] yout73;
output signed [15:0] yout74;
output signed [15:0] yout75;
output signed [15:0] yout76;
output signed [15:0] yout77;
output signed [15:0] yout78;
output signed [15:0] yout79;
output signed [15:0] yout80;
output signed [15:0] yout81;
output signed [15:0] yout82;
output signed [15:0] yout83;
output signed [15:0] yout84;
output signed [15:0] yout85;
output signed [15:0] yout86;
output signed [15:0] yout87;
output signed [15:0] yout88;
output signed [15:0] yout89;
output signed [15:0] yout90;
output signed [15:0] yout91;
output signed [15:0] yout92;
output signed [15:0] yout93;
output signed [15:0] yout94;
output signed [15:0] yout95;
output signed [15:0] yout96;
output signed [15:0] yout97;
output signed [15:0] yout98;
output signed [15:0] yout99;
output signed [15:0] yout100;
output signed [15:0] yout101;
output signed [15:0] yout102;
output signed [15:0] yout103;
output signed [15:0] yout104;
output signed [15:0] yout105;
output signed [15:0] yout106;
output signed [15:0] yout107;
output signed [15:0] yout108;
output signed [15:0] yout109;
output signed [15:0] yout110;
output signed [15:0] yout111;
output signed [15:0] yout112;
output signed [15:0] yout113;
output signed [15:0] yout114;
output signed [15:0] yout115;
output signed [15:0] yout116;
output signed [15:0] yout117;
output signed [15:0] yout118;
output signed [15:0] yout119;
output signed [15:0] yout120;
output signed [15:0] yout121;
output signed [15:0] yout122;
output signed [15:0] yout123;
output signed [15:0] yout124;
output signed [15:0] yout125;
output signed [15:0] yout126;
output signed [15:0] yout127;
output signed [15:0] yout128;
output signed [15:0] yout129;
output signed [15:0] yout130;
output signed [15:0] yout131;
output signed [15:0] yout132;
output signed [15:0] yout133;
output signed [15:0] yout134;
output signed [15:0] yout135;
output signed [15:0] yout136;
output signed [15:0] yout137;
output signed [15:0] yout138;
output signed [15:0] yout139;
output signed [15:0] yout140;
output signed [15:0] yout141;
output signed [15:0] yout142;
output signed [15:0] yout143;
output signed [15:0] yout144;
output signed [15:0] yout145;
output signed [15:0] yout146;
output signed [15:0] yout147;
output signed [15:0] yout148;
output signed [15:0] yout149;
output signed [15:0] yout150;
output signed [15:0] yout151;
output signed [15:0] yout152;
output signed [15:0] yout153;
output signed [15:0] yout154;
output signed [15:0] yout155;
output signed [15:0] yout156;
output signed [15:0] yout157;
output signed [15:0] yout158;
output signed [15:0] yout159;
output signed [15:0] yout160;
output signed [15:0] yout161;
output signed [15:0] yout162;
output signed [15:0] yout163;
output signed [15:0] yout164;
output signed [15:0] yout165;
output signed [15:0] yout166;
output signed [15:0] yout167;
output signed [15:0] yout168;
output signed [15:0] yout169;
output signed [15:0] yout170;
output signed [15:0] yout171;
output signed [15:0] yout172;
output signed [15:0] yout173;
output signed [15:0] yout174;
output signed [15:0] yout175;
output signed [15:0] yout176;
output signed [15:0] yout177;
output signed [15:0] yout178;
output signed [15:0] yout179;
output signed [15:0] yout180;
output signed [15:0] yout181;
output signed [15:0] yout182;
output signed [15:0] yout183;
output signed [15:0] yout184;
output signed [15:0] yout185;
output signed [15:0] yout186;
output signed [15:0] yout187;
output signed [15:0] yout188;
output signed [15:0] yout189;
output signed [15:0] yout190;
output signed [15:0] yout191;
output signed [15:0] yout192;
output signed [15:0] yout193;
output signed [15:0] yout194;
output signed [15:0] yout195;
output signed [15:0] yout196;
output signed [15:0] yout197;
output signed [15:0] yout198;
output signed [15:0] yout199;
output signed [15:0] yout200;
output signed [15:0] yout201;
output signed [15:0] yout202;
output signed [15:0] yout203;
output signed [15:0] yout204;
output signed [15:0] yout205;
output signed [15:0] yout206;
output signed [15:0] yout207;
output signed [15:0] yout208;
output signed [15:0] yout209;
output signed [15:0] yout210;
output signed [15:0] yout211;
output signed [15:0] yout212;
output signed [15:0] yout213;
output signed [15:0] yout214;
output signed [15:0] yout215;
output signed [15:0] yout216;
output signed [15:0] yout217;
output signed [15:0] yout218;
output signed [15:0] yout219;
output signed [15:0] yout220;
output signed [15:0] yout221;
output signed [15:0] yout222;
output signed [15:0] yout223;
output signed [15:0] yout224;
output signed [15:0] yout225;
output signed [15:0] yout226;
output signed [15:0] yout227;
output signed [15:0] yout228;
output signed [15:0] yout229;
output signed [15:0] yout230;
output signed [15:0] yout231;
output signed [15:0] yout232;
output signed [15:0] yout233;
output signed [15:0] yout234;
output signed [15:0] yout235;
output signed [15:0] yout236;
output signed [15:0] yout237;
output signed [15:0] yout238;
output signed [15:0] yout239;
output signed [15:0] yout240;
output signed [15:0] yout241;
output signed [15:0] yout242;
output signed [15:0] yout243;
output signed [15:0] yout244;
output signed [15:0] yout245;
output signed [15:0] yout246;
output signed [15:0] yout247;
output signed [15:0] yout248;
output signed [15:0] yout249;
output signed [15:0] yout250;
output signed [15:0] yout251;
output signed [15:0] yout252;
output signed [15:0] yout253;
output signed [15:0] yout254;
output signed [15:0] yout255;
output signed [15:0] yout256;
    
    
ifft ifft1(
xin1,xin2,xin3,xin4,xin5,xin6,xin7,xin8,xin9,xin10,xin11,xin12,xin13,xin14,xin15,xin16,
yin1,yin2,yin3,yin4,yin5,yin6,yin7,yin8,yin9,yin10,yin11,yin12,yin13,yin14,yin15,yin16,
clock,
xout1,xout2,xout3,xout4,xout5,xout6,xout7,xout8,xout9,xout10,xout11,xout12,xout13,xout14,xout15,xout16,
yout1,yout2,yout3,yout4,yout5,yout6,yout7,yout8,yout9,yout10,yout11,yout12,yout13,yout14,yout15,yout16
);

ifft ifft2(
xin17,xin18,xin19,xin20,xin21,xin22,xin23,xin24,xin25,xin26,xin27,xin28,xin29,xin30,xin31,xin32,
yin17,yin18,yin19,yin20,yin21,yin22,yin23,yin24,yin25,yin26,yin27,yin28,yin29,yin30,yin31,yin32,
clock,
xout17,xout18,xout19,xout20,xout21,xout22,xout23,xout24,xout25,xout26,xout27,xout28,xout29,xout30,xout31,xout32,
yout17,yout18,yout19,yout20,yout21,yout22,yout23,yout24,yout25,yout26,yout27,yout28,yout29,yout30,yout31,yout32
);

ifft ifft3(
xin33,xin34,xin35,xin36,xin37,xin38,xin39,xin40,xin41,xin42,xin43,xin44,xin45,xin46,xin47,xin48,
yin33,yin34,yin35,yin36,yin37,yin38,yin39,yin40,yin41,yin42,yin43,yin44,yin45,yin46,yin47,yin48,
clock,
xout33,xout34,xout35,xout36,xout37,xout38,xout39,xout40,xout41,xout42,xout43,xout44,xout45,xout46,xout47,xout48,
yout33,yout34,yout35,yout36,yout37,yout38,yout39,yout40,yout41,yout42,yout43,yout44,yout45,yout46,yout47,yout48
);

ifft ifft4(
xin49,xin50,xin51,xin52,xin53,xin54,xin55,xin56,xin57,xin58,xin59,xin60,xin61,xin62,xin63,xin64,
yin49,yin50,yin51,yin52,yin53,yin54,yin55,yin56,yin57,yin58,yin59,yin60,yin61,yin62,yin63,yin64,
clock,
xout49,xout50,xout51,xout52,xout53,xout54,xout55,xout56,xout57,xout58,xout59,xout60,xout61,xout62,xout63,xout64,
yout49,yout50,yout51,yout52,yout53,yout54,yout55,yout56,yout57,yout58,yout59,yout60,yout61,yout62,yout63,yout64
);

ifft ifft5(
xin65,xin66,xin67,xin68,xin69,xin70,xin71,xin72,xin73,xin74,xin75,xin76,xin77,xin78,xin79,xin80,
yin65,yin66,yin67,yin68,yin69,yin70,yin71,yin72,yin73,yin74,yin75,yin76,yin77,yin78,yin79,yin80,
clock,
xout65,xout66,xout67,xout68,xout69,xout70,xout71,xout72,xout73,xout74,xout75,xout76,xout77,xout78,xout79,xout80,
yout65,yout66,yout67,yout68,yout69,yout70,yout71,yout72,yout73,yout74,yout75,yout76,yout77,yout78,yout79,yout80
);

ifft ifft6(
xin81,xin82,xin83,xin84,xin85,xin86,xin87,xin88,xin89,xin90,xin91,xin92,xin93,xin94,xin95,xin96,
yin81,yin82,yin83,yin84,yin85,yin86,yin87,yin88,yin89,yin90,yin91,yin92,yin93,yin94,yin95,yin96,
clock,
xout81,xout82,xout83,xout84,xout85,xout86,xout87,xout88,xout89,xout90,xout91,xout92,xout93,xout94,xout95,xout96,
yout81,yout82,yout83,yout84,yout85,yout86,yout87,yout88,yout89,yout90,yout91,yout92,yout93,yout94,yout95,yout96
);

ifft ifft7(
xin97,xin98,xin99,xin100,xin101,xin102,xin103,xin104,xin105,xin106,xin107,xin108,xin109,xin110,xin111,xin112,
yin97,yin98,yin99,yin100,yin101,yin102,yin103,yin104,yin105,yin106,yin107,yin108,yin109,yin110,yin111,yin112,
clock,
xout97,xout98,xout99,xout100,xout101,xout102,xout103,xout104,xout105,xout106,xout107,xout108,xout109,xout110,xout111,xout112,
yout97,yout98,yout99,yout100,yout101,yout102,yout103,yout104,yout105,yout106,yout107,yout108,yout109,yout110,yout111,yout112
);

ifft ifft8(
xin113,xin114,xin115,xin116,xin117,xin118,xin119,xin120,xin121,xin122,xin123,xin124,xin125,xin126,xin127,xin128,
yin113,yin114,yin115,yin116,yin117,yin118,yin119,yin120,yin121,yin122,yin123,yin124,yin125,yin126,yin127,yin128,
clock,
xout113,xout114,xout115,xout116,xout117,xout118,xout119,xout120,xout121,xout122,xout123,xout124,xout125,xout126,xout127,xout128,
yout113,yout114,yout115,yout116,yout117,yout118,yout119,yout120,yout121,yout122,yout123,yout124,yout125,yout126,yout127,yout128
);

ifft ifft9(
xin129,xin130,xin131,xin132,xin133,xin134,xin135,xin136,xin137,xin138,xin139,xin140,xin141,xin142,xin143,xin144,
yin129,yin130,yin131,yin132,yin133,yin134,yin135,yin136,yin137,yin138,yin139,yin140,yin141,yin142,yin143,yin144,
clock,
xout129,xout130,xout131,xout132,xout133,xout134,xout135,xout136,xout137,xout138,xout139,xout140,xout141,xout142,xout143,xout144,
yout129,yout130,yout131,yout132,yout133,yout134,yout135,yout136,yout137,yout138,yout139,yout140,yout141,yout142,yout143,yout144
);

ifft ifft10(
xin145,xin146,xin147,xin148,xin149,xin150,xin151,xin152,xin153,xin154,xin155,xin156,xin157,xin158,xin159,xin160,
yin145,yin146,yin147,yin148,yin149,yin150,yin151,yin152,yin153,yin154,yin155,yin156,yin157,yin158,yin159,yin160,
clock,
xout145,xout146,xout147,xout148,xout149,xout150,xout151,xout152,xout153,xout154,xout155,xout156,xout157,xout158,xout159,xout160,
yout145,yout146,yout147,yout148,yout149,yout150,yout151,yout152,yout153,yout154,yout155,yout156,yout157,yout158,yout159,yout160
);

ifft ifft11(
xin161,xin162,xin163,xin164,xin165,xin166,xin167,xin168,xin169,xin170,xin171,xin172,xin173,xin174,xin175,xin176,
yin161,yin162,yin163,yin164,yin165,yin166,yin167,yin168,yin169,yin170,yin171,yin172,yin173,yin174,yin175,yin176,
clock,
xout161,xout162,xout163,xout164,xout165,xout166,xout167,xout168,xout169,xout170,xout171,xout172,xout173,xout174,xout175,xout176,
yout161,yout162,yout163,yout164,yout165,yout166,yout167,yout168,yout169,yout170,yout171,yout172,yout173,yout174,yout175,yout176
);

ifft ifft12(
xin177,xin178,xin179,xin180,xin181,xin182,xin183,xin184,xin185,xin186,xin187,xin188,xin189,xin190,xin191,xin192,
yin177,yin178,yin179,yin180,yin181,yin182,yin183,yin184,yin185,yin186,yin187,yin188,yin189,yin190,yin191,yin192,
clock,
xout177,xout178,xout179,xout180,xout181,xout182,xout183,xout184,xout185,xout186,xout187,xout188,xout189,xout190,xout191,xout192,
yout177,yout178,yout179,yout180,yout181,yout182,yout183,yout184,yout185,yout186,yout187,yout188,yout189,yout190,yout191,yout192
);

ifft ifft13(
xin193,xin194,xin195,xin196,xin197,xin198,xin199,xin200,xin201,xin202,xin203,xin204,xin205,xin206,xin207,xin208,
yin193,yin194,yin195,yin196,yin197,yin198,yin199,yin200,yin201,yin202,yin203,yin204,yin205,yin206,yin207,yin208,
clock,
xout193,xout194,xout195,xout196,xout197,xout198,xout199,xout200,xout201,xout202,xout203,xout204,xout205,xout206,xout207,xout208,
yout193,yout194,yout195,yout196,yout197,yout198,yout199,yout200,yout201,yout202,yout203,yout204,yout205,yout206,yout207,yout208
);

ifft ifft14(
xin209,xin210,xin211,xin212,xin213,xin214,xin215,xin216,xin217,xin218,xin219,xin220,xin221,xin222,xin223,xin224,
yin209,yin210,yin211,yin212,yin213,yin214,yin215,yin216,yin217,yin218,yin219,yin220,yin221,yin222,yin223,yin224,
clock,
xout209,xout210,xout211,xout212,xout213,xout214,xout215,xout216,xout217,xout218,xout219,xout220,xout221,xout222,xout223,xout224,
yout209,yout210,yout211,yout212,yout213,yout214,yout215,yout216,yout217,yout218,yout219,yout220,yout221,yout222,yout223,yout224
);

ifft ifft15(
xin225,xin226,xin227,xin228,xin229,xin230,xin231,xin232,xin233,xin234,xin235,xin236,xin237,xin238,xin239,xin240,
yin225,yin226,yin227,yin228,yin229,yin230,yin231,yin232,yin233,yin234,yin235,yin236,yin237,yin238,yin239,yin240,
clock,
xout225,xout226,xout227,xout228,xout229,xout230,xout231,xout232,xout233,xout234,xout235,xout236,xout237,xout238,xout239,xout240,
yout225,yout226,yout227,yout228,yout229,yout230,yout231,yout232,yout233,yout234,yout235,yout236,yout237,yout238,yout239,yout240
);

ifft ifft16(
xin241,xin242,xin243,xin244,xin245,xin246,xin247,xin248,xin249,xin250,xin251,xin252,xin253,xin254,xin255,xin256,
yin241,yin242,yin243,yin244,yin245,yin246,yin247,yin248,yin249,yin250,yin251,yin252,yin253,yin254,yin255,yin256,
clock,
xout241,xout242,xout243,xout244,xout245,xout246,xout247,xout248,xout249,xout250,xout251,xout252,xout253,xout254,xout255,xout256,
yout241,yout242,yout243,yout244,yout245,yout246,yout247,yout248,yout249,yout250,yout251,yout252,yout253,yout254,yout255,yout256
);

endmodule
