`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.08.2023 23:59:17
// Design Name: 
// Module Name: otfs_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module otfs_tb;

reg [15:0] xin1 =0;
reg [15:0] xin2 =0;
reg [15:0] xin3 =0;
reg [15:0] xin4 =0;
reg [15:0] xin5 =0;
reg [15:0] xin6 =0;
reg [15:0] xin7 =0;
reg [15:0] xin8 =0;
reg [15:0] xin9 =0;
reg [15:0] xin10 =0;
reg [15:0] xin11 =0;
reg [15:0] xin12 =0;
reg [15:0] xin13 =0;
reg [15:0] xin14 =0;
reg [15:0] xin15 =0;
reg [15:0] xin16 =0;
reg [15:0] xin17 =0;
reg [15:0] xin18 =0;
reg [15:0] xin19 =0;
reg [15:0] xin20 =0;
reg [15:0] xin21 =0;
reg [15:0] xin22 =0;
reg [15:0] xin23 =0;
reg [15:0] xin24 =0;
reg [15:0] xin25 =0;
reg [15:0] xin26 =0;
reg [15:0] xin27 =0;
reg [15:0] xin28 =0;
reg [15:0] xin29 =0;
reg [15:0] xin30 =0;
reg [15:0] xin31 =0;
reg [15:0] xin32 =0;
reg [15:0] xin33 =0;
reg [15:0] xin34 =0;
reg [15:0] xin35 =0;
reg [15:0] xin36 =0;
reg [15:0] xin37 =0;
reg [15:0] xin38 =0;
reg [15:0] xin39 =0;
reg [15:0] xin40 =0;
reg [15:0] xin41 =0;
reg [15:0] xin42 =0;
reg [15:0] xin43 =0;
reg [15:0] xin44 =0;
reg [15:0] xin45 =0;
reg [15:0] xin46 =0;
reg [15:0] xin47 =0;
reg [15:0] xin48 =0;
reg [15:0] xin49 =0;
reg [15:0] xin50 =0;
reg [15:0] xin51 =0;
reg [15:0] xin52 =0;
reg [15:0] xin53 =0;
reg [15:0] xin54 =0;
reg [15:0] xin55 =0;
reg [15:0] xin56 =0;
reg [15:0] xin57 =0;
reg [15:0] xin58 =0;
reg [15:0] xin59 =0;
reg [15:0] xin60 =0;
reg [15:0] xin61 =0;
reg [15:0] xin62 =0;
reg [15:0] xin63 =0;
reg [15:0] xin64 =0;
reg [15:0] xin65 =0;
reg [15:0] xin66 =0;
reg [15:0] xin67 =0;
reg [15:0] xin68 =0;
reg [15:0] xin69 =0;
reg [15:0] xin70 =0;
reg [15:0] xin71 =0;
reg [15:0] xin72 =0;
reg [15:0] xin73 =0;
reg [15:0] xin74 =0;
reg [15:0] xin75 =0;
reg [15:0] xin76 =0;
reg [15:0] xin77 =0;
reg [15:0] xin78 =0;
reg [15:0] xin79 =0;
reg [15:0] xin80 =0;
reg [15:0] xin81 =0;
reg [15:0] xin82 =0;
reg [15:0] xin83 =0;
reg [15:0] xin84 =0;
reg [15:0] xin85 =0;
reg [15:0] xin86 =0;
reg [15:0] xin87 =0;
reg [15:0] xin88 =0;
reg [15:0] xin89 =0;
reg [15:0] xin90 =0;
reg [15:0] xin91 =0;
reg [15:0] xin92 =0;
reg [15:0] xin93 =0;
reg [15:0] xin94 =0;
reg [15:0] xin95 =0;
reg [15:0] xin96 =0;
reg [15:0] xin97 =0;
reg [15:0] xin98 =0;
reg [15:0] xin99 =0;
reg [15:0] xin100 =0;
reg [15:0] xin101 =0;
reg [15:0] xin102 =0;
reg [15:0] xin103 =0;
reg [15:0] xin104 =0;
reg [15:0] xin105 =0;
reg [15:0] xin106 =0;
reg [15:0] xin107 =0;
reg [15:0] xin108 =0;
reg [15:0] xin109 =0;
reg [15:0] xin110 =0;
reg [15:0] xin111 =0;
reg [15:0] xin112 =0;
reg [15:0] xin113 =0;
reg [15:0] xin114 =0;
reg [15:0] xin115 =0;
reg [15:0] xin116 =0;
reg [15:0] xin117 =0;
reg [15:0] xin118 =0;
reg [15:0] xin119 =0;
reg [15:0] xin120 =0;
reg [15:0] xin121 =0;
reg [15:0] xin122 =0;
reg [15:0] xin123 =0;
reg [15:0] xin124 =0;
reg [15:0] xin125 =0;
reg [15:0] xin126 =0;
reg [15:0] xin127 =0;
reg [15:0] xin128 =0;
reg [15:0] xin129 =0;
reg [15:0] xin130 =0;
reg [15:0] xin131 =0;
reg [15:0] xin132 =0;
reg [15:0] xin133 =0;
reg [15:0] xin134 =0;
reg [15:0] xin135 =0;
reg [15:0] xin136 =0;
reg [15:0] xin137 =0;
reg [15:0] xin138 =0;
reg [15:0] xin139 =0;
reg [15:0] xin140 =0;
reg [15:0] xin141 =0;
reg [15:0] xin142 =0;
reg [15:0] xin143 =0;
reg [15:0] xin144 =0;
reg [15:0] xin145 =0;
reg [15:0] xin146 =0;
reg [15:0] xin147 =0;
reg [15:0] xin148 =0;
reg [15:0] xin149 =0;
reg [15:0] xin150 =0;
reg [15:0] xin151 =0;
reg [15:0] xin152 =0;
reg [15:0] xin153 =0;
reg [15:0] xin154 =0;
reg [15:0] xin155 =0;
reg [15:0] xin156 =0;
reg [15:0] xin157 =0;
reg [15:0] xin158 =0;
reg [15:0] xin159 =0;
reg [15:0] xin160 =0;
reg [15:0] xin161 =0;
reg [15:0] xin162 =0;
reg [15:0] xin163 =0;
reg [15:0] xin164 =0;
reg [15:0] xin165 =0;
reg [15:0] xin166 =0;
reg [15:0] xin167 =0;
reg [15:0] xin168 =0;
reg [15:0] xin169 =0;
reg [15:0] xin170 =0;
reg [15:0] xin171 =0;
reg [15:0] xin172 =0;
reg [15:0] xin173 =0;
reg [15:0] xin174 =0;
reg [15:0] xin175 =0;
reg [15:0] xin176 =0;
reg [15:0] xin177 =0;
reg [15:0] xin178 =0;
reg [15:0] xin179 =0;
reg [15:0] xin180 =0;
reg [15:0] xin181 =0;
reg [15:0] xin182 =0;
reg [15:0] xin183 =0;
reg [15:0] xin184 =0;
reg [15:0] xin185 =0;
reg [15:0] xin186 =0;
reg [15:0] xin187 =0;
reg [15:0] xin188 =0;
reg [15:0] xin189 =0;
reg [15:0] xin190 =0;
reg [15:0] xin191 =0;
reg [15:0] xin192 =0;
reg [15:0] xin193 =0;
reg [15:0] xin194 =0;
reg [15:0] xin195 =0;
reg [15:0] xin196 =0;
reg [15:0] xin197 =0;
reg [15:0] xin198 =0;
reg [15:0] xin199 =0;
reg [15:0] xin200 =0;
reg [15:0] xin201 =0;
reg [15:0] xin202 =0;
reg [15:0] xin203 =0;
reg [15:0] xin204 =0;
reg [15:0] xin205 =0;
reg [15:0] xin206 =0;
reg [15:0] xin207 =0;
reg [15:0] xin208 =0;
reg [15:0] xin209 =0;
reg [15:0] xin210 =0;
reg [15:0] xin211 =0;
reg [15:0] xin212 =0;
reg [15:0] xin213 =0;
reg [15:0] xin214 =0;
reg [15:0] xin215 =0;
reg [15:0] xin216 =0;
reg [15:0] xin217 =0;
reg [15:0] xin218 =0;
reg [15:0] xin219 =0;
reg [15:0] xin220 =0;
reg [15:0] xin221 =0;
reg [15:0] xin222 =0;
reg [15:0] xin223 =0;
reg [15:0] xin224 =0;
reg [15:0] xin225 =0;
reg [15:0] xin226 =0;
reg [15:0] xin227 =0;
reg [15:0] xin228 =0;
reg [15:0] xin229 =0;
reg [15:0] xin230 =0;
reg [15:0] xin231 =0;
reg [15:0] xin232 =0;
reg [15:0] xin233 =0;
reg [15:0] xin234 =0;
reg [15:0] xin235 =0;
reg [15:0] xin236 =0;
reg [15:0] xin237 =0;
reg [15:0] xin238 =0;
reg [15:0] xin239 =0;
reg [15:0] xin240 =0;
reg [15:0] xin241 =0;
reg [15:0] xin242 =0;
reg [15:0] xin243 =0;
reg [15:0] xin244 =0;
reg [15:0] xin245 =0;
reg [15:0] xin246 =0;
reg [15:0] xin247 =0;
reg [15:0] xin248 =0;
reg [15:0] xin249 =0;
reg [15:0] xin250 =0;
reg [15:0] xin251 =0;
reg [15:0] xin252 =0;
reg [15:0] xin253 =0;
reg [15:0] xin254 =0;
reg [15:0] xin255 =0;
reg [15:0] xin256 =0;

reg [15:0] yin1 =0;
reg [15:0] yin2 =0;
reg [15:0] yin3 =0;
reg [15:0] yin4 =0;
reg [15:0] yin5 =0;
reg [15:0] yin6 =0;
reg [15:0] yin7 =0;
reg [15:0] yin8 =0;
reg [15:0] yin9 =0;
reg [15:0] yin10 =0;
reg [15:0] yin11 =0;
reg [15:0] yin12 =0;
reg [15:0] yin13 =0;
reg [15:0] yin14 =0;
reg [15:0] yin15 =0;
reg [15:0] yin16 =0;
reg [15:0] yin17 =0;
reg [15:0] yin18 =0;
reg [15:0] yin19 =0;
reg [15:0] yin20 =0;
reg [15:0] yin21 =0;
reg [15:0] yin22 =0;
reg [15:0] yin23 =0;
reg [15:0] yin24 =0;
reg [15:0] yin25 =0;
reg [15:0] yin26 =0;
reg [15:0] yin27 =0;
reg [15:0] yin28 =0;
reg [15:0] yin29 =0;
reg [15:0] yin30 =0;
reg [15:0] yin31 =0;
reg [15:0] yin32 =0;
reg [15:0] yin33 =0;
reg [15:0] yin34 =0;
reg [15:0] yin35 =0;
reg [15:0] yin36 =0;
reg [15:0] yin37 =0;
reg [15:0] yin38 =0;
reg [15:0] yin39 =0;
reg [15:0] yin40 =0;
reg [15:0] yin41 =0;
reg [15:0] yin42 =0;
reg [15:0] yin43 =0;
reg [15:0] yin44 =0;
reg [15:0] yin45 =0;
reg [15:0] yin46 =0;
reg [15:0] yin47 =0;
reg [15:0] yin48 =0;
reg [15:0] yin49 =0;
reg [15:0] yin50 =0;
reg [15:0] yin51 =0;
reg [15:0] yin52 =0;
reg [15:0] yin53 =0;
reg [15:0] yin54 =0;
reg [15:0] yin55 =0;
reg [15:0] yin56 =0;
reg [15:0] yin57 =0;
reg [15:0] yin58 =0;
reg [15:0] yin59 =0;
reg [15:0] yin60 =0;
reg [15:0] yin61 =0;
reg [15:0] yin62 =0;
reg [15:0] yin63 =0;
reg [15:0] yin64 =0;
reg [15:0] yin65 =0;
reg [15:0] yin66 =0;
reg [15:0] yin67 =0;
reg [15:0] yin68 =0;
reg [15:0] yin69 =0;
reg [15:0] yin70 =0;
reg [15:0] yin71 =0;
reg [15:0] yin72 =0;
reg [15:0] yin73 =0;
reg [15:0] yin74 =0;
reg [15:0] yin75 =0;
reg [15:0] yin76 =0;
reg [15:0] yin77 =0;
reg [15:0] yin78 =0;
reg [15:0] yin79 =0;
reg [15:0] yin80 =0;
reg [15:0] yin81 =0;
reg [15:0] yin82 =0;
reg [15:0] yin83 =0;
reg [15:0] yin84 =0;
reg [15:0] yin85 =0;
reg [15:0] yin86 =0;
reg [15:0] yin87 =0;
reg [15:0] yin88 =0;
reg [15:0] yin89 =0;
reg [15:0] yin90 =0;
reg [15:0] yin91 =0;
reg [15:0] yin92 =0;
reg [15:0] yin93 =0;
reg [15:0] yin94 =0;
reg [15:0] yin95 =0;
reg [15:0] yin96 =0;
reg [15:0] yin97 =0;
reg [15:0] yin98 =0;
reg [15:0] yin99 =0;
reg [15:0] yin100 =0;
reg [15:0] yin101 =0;
reg [15:0] yin102 =0;
reg [15:0] yin103 =0;
reg [15:0] yin104 =0;
reg [15:0] yin105 =0;
reg [15:0] yin106 =0;
reg [15:0] yin107 =0;
reg [15:0] yin108 =0;
reg [15:0] yin109 =0;
reg [15:0] yin110 =0;
reg [15:0] yin111 =0;
reg [15:0] yin112 =0;
reg [15:0] yin113 =0;
reg [15:0] yin114 =0;
reg [15:0] yin115 =0;
reg [15:0] yin116 =0;
reg [15:0] yin117 =0;
reg [15:0] yin118 =0;
reg [15:0] yin119 =0;
reg [15:0] yin120 =0;
reg [15:0] yin121 =0;
reg [15:0] yin122 =0;
reg [15:0] yin123 =0;
reg [15:0] yin124 =0;
reg [15:0] yin125 =0;
reg [15:0] yin126 =0;
reg [15:0] yin127 =0;
reg [15:0] yin128 =0;
reg [15:0] yin129 =0;
reg [15:0] yin130 =0;
reg [15:0] yin131 =0;
reg [15:0] yin132 =0;
reg [15:0] yin133 =0;
reg [15:0] yin134 =0;
reg [15:0] yin135 =0;
reg [15:0] yin136 =0;
reg [15:0] yin137 =0;
reg [15:0] yin138 =0;
reg [15:0] yin139 =0;
reg [15:0] yin140 =0;
reg [15:0] yin141 =0;
reg [15:0] yin142 =0;
reg [15:0] yin143 =0;
reg [15:0] yin144 =0;
reg [15:0] yin145 =0;
reg [15:0] yin146 =0;
reg [15:0] yin147 =0;
reg [15:0] yin148 =0;
reg [15:0] yin149 =0;
reg [15:0] yin150 =0;
reg [15:0] yin151 =0;
reg [15:0] yin152 =0;
reg [15:0] yin153 =0;
reg [15:0] yin154 =0;
reg [15:0] yin155 =0;
reg [15:0] yin156 =0;
reg [15:0] yin157 =0;
reg [15:0] yin158 =0;
reg [15:0] yin159 =0;
reg [15:0] yin160 =0;
reg [15:0] yin161 =0;
reg [15:0] yin162 =0;
reg [15:0] yin163 =0;
reg [15:0] yin164 =0;
reg [15:0] yin165 =0;
reg [15:0] yin166 =0;
reg [15:0] yin167 =0;
reg [15:0] yin168 =0;
reg [15:0] yin169 =0;
reg [15:0] yin170 =0;
reg [15:0] yin171 =0;
reg [15:0] yin172 =0;
reg [15:0] yin173 =0;
reg [15:0] yin174 =0;
reg [15:0] yin175 =0;
reg [15:0] yin176 =0;
reg [15:0] yin177 =0;
reg [15:0] yin178 =0;
reg [15:0] yin179 =0;
reg [15:0] yin180 =0;
reg [15:0] yin181 =0;
reg [15:0] yin182 =0;
reg [15:0] yin183 =0;
reg [15:0] yin184 =0;
reg [15:0] yin185 =0;
reg [15:0] yin186 =0;
reg [15:0] yin187 =0;
reg [15:0] yin188 =0;
reg [15:0] yin189 =0;
reg [15:0] yin190 =0;
reg [15:0] yin191 =0;
reg [15:0] yin192 =0;
reg [15:0] yin193 =0;
reg [15:0] yin194 =0;
reg [15:0] yin195 =0;
reg [15:0] yin196 =0;
reg [15:0] yin197 =0;
reg [15:0] yin198 =0;
reg [15:0] yin199 =0;
reg [15:0] yin200 =0;
reg [15:0] yin201 =0;
reg [15:0] yin202 =0;
reg [15:0] yin203 =0;
reg [15:0] yin204 =0;
reg [15:0] yin205 =0;
reg [15:0] yin206 =0;
reg [15:0] yin207 =0;
reg [15:0] yin208 =0;
reg [15:0] yin209 =0;
reg [15:0] yin210 =0;
reg [15:0] yin211 =0;
reg [15:0] yin212 =0;
reg [15:0] yin213 =0;
reg [15:0] yin214 =0;
reg [15:0] yin215 =0;
reg [15:0] yin216 =0;
reg [15:0] yin217 =0;
reg [15:0] yin218 =0;
reg [15:0] yin219 =0;
reg [15:0] yin220 =0;
reg [15:0] yin221 =0;
reg [15:0] yin222 =0;
reg [15:0] yin223 =0;
reg [15:0] yin224 =0;
reg [15:0] yin225 =0;
reg [15:0] yin226 =0;
reg [15:0] yin227 =0;
reg [15:0] yin228 =0;
reg [15:0] yin229 =0;
reg [15:0] yin230 =0;
reg [15:0] yin231 =0;
reg [15:0] yin232 =0;
reg [15:0] yin233 =0;
reg [15:0] yin234 =0;
reg [15:0] yin235 =0;
reg [15:0] yin236 =0;
reg [15:0] yin237 =0;
reg [15:0] yin238 =0;
reg [15:0] yin239 =0;
reg [15:0] yin240 =0;
reg [15:0] yin241 =0;
reg [15:0] yin242 =0;
reg [15:0] yin243 =0;
reg [15:0] yin244 =0;
reg [15:0] yin245 =0;
reg [15:0] yin246 =0;
reg [15:0] yin247 =0;
reg [15:0] yin248 =0;
reg [15:0] yin249 =0;
reg [15:0] yin250 =0;
reg [15:0] yin251 =0;
reg [15:0] yin252 =0;
reg [15:0] yin253 =0;
reg [15:0] yin254 =0;
reg [15:0] yin255 =0;
reg [15:0] yin256 =0;

reg clock=0;

wire [15:0] xout1;
wire [15:0] xout2;
wire [15:0] xout3;
wire [15:0] xout4;
wire [15:0] xout5;
wire [15:0] xout6;
wire [15:0] xout7;
wire [15:0] xout8;
wire [15:0] xout9;
wire [15:0] xout10;
wire [15:0] xout11;
wire [15:0] xout12;
wire [15:0] xout13;
wire [15:0] xout14;
wire [15:0] xout15;
wire [15:0] xout16;
wire [15:0] xout17;
wire [15:0] xout18;
wire [15:0] xout19;
wire [15:0] xout20;
wire [15:0] xout21;
wire [15:0] xout22;
wire [15:0] xout23;
wire [15:0] xout24;
wire [15:0] xout25;
wire [15:0] xout26;
wire [15:0] xout27;
wire [15:0] xout28;
wire [15:0] xout29;
wire [15:0] xout30;
wire [15:0] xout31;
wire [15:0] xout32;
wire [15:0] xout33;
wire [15:0] xout34;
wire [15:0] xout35;
wire [15:0] xout36;
wire [15:0] xout37;
wire [15:0] xout38;
wire [15:0] xout39;
wire [15:0] xout40;
wire [15:0] xout41;
wire [15:0] xout42;
wire [15:0] xout43;
wire [15:0] xout44;
wire [15:0] xout45;
wire [15:0] xout46;
wire [15:0] xout47;
wire [15:0] xout48;
wire [15:0] xout49;
wire [15:0] xout50;
wire [15:0] xout51;
wire [15:0] xout52;
wire [15:0] xout53;
wire [15:0] xout54;
wire [15:0] xout55;
wire [15:0] xout56;
wire [15:0] xout57;
wire [15:0] xout58;
wire [15:0] xout59;
wire [15:0] xout60;
wire [15:0] xout61;
wire [15:0] xout62;
wire [15:0] xout63;
wire [15:0] xout64;
wire [15:0] xout65;
wire [15:0] xout66;
wire [15:0] xout67;
wire [15:0] xout68;
wire [15:0] xout69;
wire [15:0] xout70;
wire [15:0] xout71;
wire [15:0] xout72;
wire [15:0] xout73;
wire [15:0] xout74;
wire [15:0] xout75;
wire [15:0] xout76;
wire [15:0] xout77;
wire [15:0] xout78;
wire [15:0] xout79;
wire [15:0] xout80;
wire [15:0] xout81;
wire [15:0] xout82;
wire [15:0] xout83;
wire [15:0] xout84;
wire [15:0] xout85;
wire [15:0] xout86;
wire [15:0] xout87;
wire [15:0] xout88;
wire [15:0] xout89;
wire [15:0] xout90;
wire [15:0] xout91;
wire [15:0] xout92;
wire [15:0] xout93;
wire [15:0] xout94;
wire [15:0] xout95;
wire [15:0] xout96;
wire [15:0] xout97;
wire [15:0] xout98;
wire [15:0] xout99;
wire [15:0] xout100;
wire [15:0] xout101;
wire [15:0] xout102;
wire [15:0] xout103;
wire [15:0] xout104;
wire [15:0] xout105;
wire [15:0] xout106;
wire [15:0] xout107;
wire [15:0] xout108;
wire [15:0] xout109;
wire [15:0] xout110;
wire [15:0] xout111;
wire [15:0] xout112;
wire [15:0] xout113;
wire [15:0] xout114;
wire [15:0] xout115;
wire [15:0] xout116;
wire [15:0] xout117;
wire [15:0] xout118;
wire [15:0] xout119;
wire [15:0] xout120;
wire [15:0] xout121;
wire [15:0] xout122;
wire [15:0] xout123;
wire [15:0] xout124;
wire [15:0] xout125;
wire [15:0] xout126;
wire [15:0] xout127;
wire [15:0] xout128;
wire [15:0] xout129;
wire [15:0] xout130;
wire [15:0] xout131;
wire [15:0] xout132;
wire [15:0] xout133;
wire [15:0] xout134;
wire [15:0] xout135;
wire [15:0] xout136;
wire [15:0] xout137;
wire [15:0] xout138;
wire [15:0] xout139;
wire [15:0] xout140;
wire [15:0] xout141;
wire [15:0] xout142;
wire [15:0] xout143;
wire [15:0] xout144;
wire [15:0] xout145;
wire [15:0] xout146;
wire [15:0] xout147;
wire [15:0] xout148;
wire [15:0] xout149;
wire [15:0] xout150;
wire [15:0] xout151;
wire [15:0] xout152;
wire [15:0] xout153;
wire [15:0] xout154;
wire [15:0] xout155;
wire [15:0] xout156;
wire [15:0] xout157;
wire [15:0] xout158;
wire [15:0] xout159;
wire [15:0] xout160;
wire [15:0] xout161;
wire [15:0] xout162;
wire [15:0] xout163;
wire [15:0] xout164;
wire [15:0] xout165;
wire [15:0] xout166;
wire [15:0] xout167;
wire [15:0] xout168;
wire [15:0] xout169;
wire [15:0] xout170;
wire [15:0] xout171;
wire [15:0] xout172;
wire [15:0] xout173;
wire [15:0] xout174;
wire [15:0] xout175;
wire [15:0] xout176;
wire [15:0] xout177;
wire [15:0] xout178;
wire [15:0] xout179;
wire [15:0] xout180;
wire [15:0] xout181;
wire [15:0] xout182;
wire [15:0] xout183;
wire [15:0] xout184;
wire [15:0] xout185;
wire [15:0] xout186;
wire [15:0] xout187;
wire [15:0] xout188;
wire [15:0] xout189;
wire [15:0] xout190;
wire [15:0] xout191;
wire [15:0] xout192;
wire [15:0] xout193;
wire [15:0] xout194;
wire [15:0] xout195;
wire [15:0] xout196;
wire [15:0] xout197;
wire [15:0] xout198;
wire [15:0] xout199;
wire [15:0] xout200;
wire [15:0] xout201;
wire [15:0] xout202;
wire [15:0] xout203;
wire [15:0] xout204;
wire [15:0] xout205;
wire [15:0] xout206;
wire [15:0] xout207;
wire [15:0] xout208;
wire [15:0] xout209;
wire [15:0] xout210;
wire [15:0] xout211;
wire [15:0] xout212;
wire [15:0] xout213;
wire [15:0] xout214;
wire [15:0] xout215;
wire [15:0] xout216;
wire [15:0] xout217;
wire [15:0] xout218;
wire [15:0] xout219;
wire [15:0] xout220;
wire [15:0] xout221;
wire [15:0] xout222;
wire [15:0] xout223;
wire [15:0] xout224;
wire [15:0] xout225;
wire [15:0] xout226;
wire [15:0] xout227;
wire [15:0] xout228;
wire [15:0] xout229;
wire [15:0] xout230;
wire [15:0] xout231;
wire [15:0] xout232;
wire [15:0] xout233;
wire [15:0] xout234;
wire [15:0] xout235;
wire [15:0] xout236;
wire [15:0] xout237;
wire [15:0] xout238;
wire [15:0] xout239;
wire [15:0] xout240;
wire [15:0] xout241;
wire [15:0] xout242;
wire [15:0] xout243;
wire [15:0] xout244;
wire [15:0] xout245;
wire [15:0] xout246;
wire [15:0] xout247;
wire [15:0] xout248;
wire [15:0] xout249;
wire [15:0] xout250;
wire [15:0] xout251;
wire [15:0] xout252;
wire [15:0] xout253;
wire [15:0] xout254;
wire [15:0] xout255;
wire [15:0] xout256;

wire [15:0] yout1;
wire [15:0] yout2;
wire [15:0] yout3;
wire [15:0] yout4;
wire [15:0] yout5;
wire [15:0] yout6;
wire [15:0] yout7;
wire [15:0] yout8;
wire [15:0] yout9;
wire [15:0] yout10;
wire [15:0] yout11;
wire [15:0] yout12;
wire [15:0] yout13;
wire [15:0] yout14;
wire [15:0] yout15;
wire [15:0] yout16;
wire [15:0] yout17;
wire [15:0] yout18;
wire [15:0] yout19;
wire [15:0] yout20;
wire [15:0] yout21;
wire [15:0] yout22;
wire [15:0] yout23;
wire [15:0] yout24;
wire [15:0] yout25;
wire [15:0] yout26;
wire [15:0] yout27;
wire [15:0] yout28;
wire [15:0] yout29;
wire [15:0] yout30;
wire [15:0] yout31;
wire [15:0] yout32;
wire [15:0] yout33;
wire [15:0] yout34;
wire [15:0] yout35;
wire [15:0] yout36;
wire [15:0] yout37;
wire [15:0] yout38;
wire [15:0] yout39;
wire [15:0] yout40;
wire [15:0] yout41;
wire [15:0] yout42;
wire [15:0] yout43;
wire [15:0] yout44;
wire [15:0] yout45;
wire [15:0] yout46;
wire [15:0] yout47;
wire [15:0] yout48;
wire [15:0] yout49;
wire [15:0] yout50;
wire [15:0] yout51;
wire [15:0] yout52;
wire [15:0] yout53;
wire [15:0] yout54;
wire [15:0] yout55;
wire [15:0] yout56;
wire [15:0] yout57;
wire [15:0] yout58;
wire [15:0] yout59;
wire [15:0] yout60;
wire [15:0] yout61;
wire [15:0] yout62;
wire [15:0] yout63;
wire [15:0] yout64;
wire [15:0] yout65;
wire [15:0] yout66;
wire [15:0] yout67;
wire [15:0] yout68;
wire [15:0] yout69;
wire [15:0] yout70;
wire [15:0] yout71;
wire [15:0] yout72;
wire [15:0] yout73;
wire [15:0] yout74;
wire [15:0] yout75;
wire [15:0] yout76;
wire [15:0] yout77;
wire [15:0] yout78;
wire [15:0] yout79;
wire [15:0] yout80;
wire [15:0] yout81;
wire [15:0] yout82;
wire [15:0] yout83;
wire [15:0] yout84;
wire [15:0] yout85;
wire [15:0] yout86;
wire [15:0] yout87;
wire [15:0] yout88;
wire [15:0] yout89;
wire [15:0] yout90;
wire [15:0] yout91;
wire [15:0] yout92;
wire [15:0] yout93;
wire [15:0] yout94;
wire [15:0] yout95;
wire [15:0] yout96;
wire [15:0] yout97;
wire [15:0] yout98;
wire [15:0] yout99;
wire [15:0] yout100;
wire [15:0] yout101;
wire [15:0] yout102;
wire [15:0] yout103;
wire [15:0] yout104;
wire [15:0] yout105;
wire [15:0] yout106;
wire [15:0] yout107;
wire [15:0] yout108;
wire [15:0] yout109;
wire [15:0] yout110;
wire [15:0] yout111;
wire [15:0] yout112;
wire [15:0] yout113;
wire [15:0] yout114;
wire [15:0] yout115;
wire [15:0] yout116;
wire [15:0] yout117;
wire [15:0] yout118;
wire [15:0] yout119;
wire [15:0] yout120;
wire [15:0] yout121;
wire [15:0] yout122;
wire [15:0] yout123;
wire [15:0] yout124;
wire [15:0] yout125;
wire [15:0] yout126;
wire [15:0] yout127;
wire [15:0] yout128;
wire [15:0] yout129;
wire [15:0] yout130;
wire [15:0] yout131;
wire [15:0] yout132;
wire [15:0] yout133;
wire [15:0] yout134;
wire [15:0] yout135;
wire [15:0] yout136;
wire [15:0] yout137;
wire [15:0] yout138;
wire [15:0] yout139;
wire [15:0] yout140;
wire [15:0] yout141;
wire [15:0] yout142;
wire [15:0] yout143;
wire [15:0] yout144;
wire [15:0] yout145;
wire [15:0] yout146;
wire [15:0] yout147;
wire [15:0] yout148;
wire [15:0] yout149;
wire [15:0] yout150;
wire [15:0] yout151;
wire [15:0] yout152;
wire [15:0] yout153;
wire [15:0] yout154;
wire [15:0] yout155;
wire [15:0] yout156;
wire [15:0] yout157;
wire [15:0] yout158;
wire [15:0] yout159;
wire [15:0] yout160;
wire [15:0] yout161;
wire [15:0] yout162;
wire [15:0] yout163;
wire [15:0] yout164;
wire [15:0] yout165;
wire [15:0] yout166;
wire [15:0] yout167;
wire [15:0] yout168;
wire [15:0] yout169;
wire [15:0] yout170;
wire [15:0] yout171;
wire [15:0] yout172;
wire [15:0] yout173;
wire [15:0] yout174;
wire [15:0] yout175;
wire [15:0] yout176;
wire [15:0] yout177;
wire [15:0] yout178;
wire [15:0] yout179;
wire [15:0] yout180;
wire [15:0] yout181;
wire [15:0] yout182;
wire [15:0] yout183;
wire [15:0] yout184;
wire [15:0] yout185;
wire [15:0] yout186;
wire [15:0] yout187;
wire [15:0] yout188;
wire [15:0] yout189;
wire [15:0] yout190;
wire [15:0] yout191;
wire [15:0] yout192;
wire [15:0] yout193;
wire [15:0] yout194;
wire [15:0] yout195;
wire [15:0] yout196;
wire [15:0] yout197;
wire [15:0] yout198;
wire [15:0] yout199;
wire [15:0] yout200;
wire [15:0] yout201;
wire [15:0] yout202;
wire [15:0] yout203;
wire [15:0] yout204;
wire [15:0] yout205;
wire [15:0] yout206;
wire [15:0] yout207;
wire [15:0] yout208;
wire [15:0] yout209;
wire [15:0] yout210;
wire [15:0] yout211;
wire [15:0] yout212;
wire [15:0] yout213;
wire [15:0] yout214;
wire [15:0] yout215;
wire [15:0] yout216;
wire [15:0] yout217;
wire [15:0] yout218;
wire [15:0] yout219;
wire [15:0] yout220;
wire [15:0] yout221;
wire [15:0] yout222;
wire [15:0] yout223;
wire [15:0] yout224;
wire [15:0] yout225;
wire [15:0] yout226;
wire [15:0] yout227;
wire [15:0] yout228;
wire [15:0] yout229;
wire [15:0] yout230;
wire [15:0] yout231;
wire [15:0] yout232;
wire [15:0] yout233;
wire [15:0] yout234;
wire [15:0] yout235;
wire [15:0] yout236;
wire [15:0] yout237;
wire [15:0] yout238;
wire [15:0] yout239;
wire [15:0] yout240;
wire [15:0] yout241;
wire [15:0] yout242;
wire [15:0] yout243;
wire [15:0] yout244;
wire [15:0] yout245;
wire [15:0] yout246;
wire [15:0] yout247;
wire [15:0] yout248;
wire [15:0] yout249;
wire [15:0] yout250;
wire [15:0] yout251;
wire [15:0] yout252;
wire [15:0] yout253;
wire [15:0] yout254;
wire [15:0] yout255;
wire [15:0] yout256;

otfs dut(       xin1, xin2, xin3, xin4, xin5, xin6, xin7, xin8, xin9, xin10, xin11, xin12, xin13, xin14, xin15, xin16, xin17, xin18, xin19, xin20, xin21, xin22, xin23, xin24, xin25, xin26, xin27, xin28, xin29, xin30, xin31, xin32, xin33, xin34, xin35, xin36, xin37, xin38, xin39, xin40, xin41, xin42, xin43, xin44, xin45, xin46, xin47, xin48, xin49, xin50, xin51, xin52, xin53, xin54, xin55, xin56, xin57, xin58, xin59, xin60, xin61, xin62, xin63, xin64, xin65, xin66, xin67, xin68, xin69, xin70, xin71, xin72, xin73, xin74, xin75, xin76, xin77, xin78, xin79, xin80, xin81, xin82, xin83, xin84, xin85, xin86, xin87, xin88, xin89, xin90, xin91, xin92, xin93, xin94, xin95, xin96, xin97, xin98, xin99, xin100, xin101, xin102, xin103, xin104, xin105, xin106, xin107, xin108, xin109, xin110, xin111, xin112, xin113, xin114, xin115, xin116, xin117, xin118, xin119, xin120, xin121, xin122, xin123, xin124, xin125, xin126, xin127, xin128, xin129, xin130, xin131, xin132, xin133, xin134, xin135, xin136, xin137, xin138, xin139, xin140, xin141, xin142, xin143, xin144, xin145, xin146, xin147, xin148, xin149, xin150, xin151, xin152, xin153, xin154, xin155, xin156, xin157, xin158, xin159, xin160, xin161, xin162, xin163, xin164, xin165, xin166, xin167, xin168, xin169, xin170, xin171, xin172, xin173, xin174, xin175, xin176, xin177, xin178, xin179, xin180, xin181, xin182, xin183, xin184, xin185, xin186, xin187, xin188, xin189, xin190, xin191, xin192, xin193, xin194, xin195, xin196, xin197, xin198, xin199, xin200, xin201, xin202, xin203, xin204, xin205, xin206, xin207, xin208, xin209, xin210, xin211, xin212, xin213, xin214, xin215, xin216, xin217, xin218, xin219, xin220, xin221, xin222, xin223, xin224, xin225, xin226, xin227, xin228, xin229, xin230, xin231, xin232, xin233, xin234, xin235, xin236, xin237, xin238, xin239, xin240, xin241, xin242, xin243, xin244, xin245, xin246, xin247, xin248, xin249, xin250, xin251, xin252, xin253, xin254, xin255, xin256,
                yin1, yin2, yin3, yin4, yin5, yin6, yin7, yin8, yin9, yin10, yin11, yin12, yin13, yin14, yin15, yin16, yin17, yin18, yin19, yin20, yin21, yin22, yin23, yin24, yin25, yin26, yin27, yin28, yin29, yin30, yin31, yin32, yin33, yin34, yin35, yin36, yin37, yin38, yin39, yin40, yin41, yin42, yin43, yin44, yin45, yin46, yin47, yin48, yin49, yin50, yin51, yin52, yin53, yin54, yin55, yin56, yin57, yin58, yin59, yin60, yin61, yin62, yin63, yin64, yin65, yin66, yin67, yin68, yin69, yin70, yin71, yin72, yin73, yin74, yin75, yin76, yin77, yin78, yin79, yin80, yin81, yin82, yin83, yin84, yin85, yin86, yin87, yin88, yin89, yin90, yin91, yin92, yin93, yin94, yin95, yin96, yin97, yin98, yin99, yin100, yin101, yin102, yin103, yin104, yin105, yin106, yin107, yin108, yin109, yin110, yin111, yin112, yin113, yin114, yin115, yin116, yin117, yin118, yin119, yin120, yin121, yin122, yin123, yin124, yin125, yin126, yin127, yin128, yin129, yin130, yin131, yin132, yin133, yin134, yin135, yin136, yin137, yin138, yin139, yin140, yin141, yin142, yin143, yin144, yin145, yin146, yin147, yin148, yin149, yin150, yin151, yin152, yin153, yin154, yin155, yin156, yin157, yin158, yin159, yin160, yin161, yin162, yin163, yin164, yin165, yin166, yin167, yin168, yin169, yin170, yin171, yin172, yin173, yin174, yin175, yin176, yin177, yin178, yin179, yin180, yin181, yin182, yin183, yin184, yin185, yin186, yin187, yin188, yin189, yin190, yin191, yin192, yin193, yin194, yin195, yin196, yin197, yin198, yin199, yin200, yin201, yin202, yin203, yin204, yin205, yin206, yin207, yin208, yin209, yin210, yin211, yin212, yin213, yin214, yin215, yin216, yin217, yin218, yin219, yin220, yin221, yin222, yin223, yin224, yin225, yin226, yin227, yin228, yin229, yin230, yin231, yin232, yin233, yin234, yin235, yin236, yin237, yin238, yin239, yin240, yin241, yin242, yin243, yin244, yin245, yin246, yin247, yin248, yin249, yin250, yin251, yin252, yin253, yin254, yin255, yin256,
                clock,
                xout1, xout2, xout3, xout4, xout5, xout6, xout7, xout8, xout9, xout10, xout11, xout12, xout13, xout14, xout15, xout16, xout17, xout18, xout19, xout20, xout21, xout22, xout23, xout24, xout25, xout26, xout27, xout28, xout29, xout30, xout31, xout32, xout33, xout34, xout35, xout36, xout37, xout38, xout39, xout40, xout41, xout42, xout43, xout44, xout45, xout46, xout47, xout48, xout49, xout50, xout51, xout52, xout53, xout54, xout55, xout56, xout57, xout58, xout59, xout60, xout61, xout62, xout63, xout64, xout65, xout66, xout67, xout68, xout69, xout70, xout71, xout72, xout73, xout74, xout75, xout76, xout77, xout78, xout79, xout80, xout81, xout82, xout83, xout84, xout85, xout86, xout87, xout88, xout89, xout90, xout91, xout92, xout93, xout94, xout95, xout96, xout97, xout98, xout99, xout100, xout101, xout102, xout103, xout104, xout105, xout106, xout107, xout108, xout109, xout110, xout111, xout112, xout113, xout114, xout115, xout116, xout117, xout118, xout119, xout120, xout121, xout122, xout123, xout124, xout125, xout126, xout127, xout128, xout129, xout130, xout131, xout132, xout133, xout134, xout135, xout136, xout137, xout138, xout139, xout140, xout141, xout142, xout143, xout144, xout145, xout146, xout147, xout148, xout149, xout150, xout151, xout152, xout153, xout154, xout155, xout156, xout157, xout158, xout159, xout160, xout161, xout162, xout163, xout164, xout165, xout166, xout167, xout168, xout169, xout170, xout171, xout172, xout173, xout174, xout175, xout176, xout177, xout178, xout179, xout180, xout181, xout182, xout183, xout184, xout185, xout186, xout187, xout188, xout189, xout190, xout191, xout192, xout193, xout194, xout195, xout196, xout197, xout198, xout199, xout200, xout201, xout202, xout203, xout204, xout205, xout206, xout207, xout208, xout209, xout210, xout211, xout212, xout213, xout214, xout215, xout216, xout217, xout218, xout219, xout220, xout221, xout222, xout223, xout224, xout225, xout226, xout227, xout228, xout229, xout230, xout231, xout232, xout233, xout234, xout235, xout236, xout237, xout238, xout239, xout240, xout241, xout242, xout243, xout244, xout245, xout246, xout247, xout248, xout249, xout250, xout251, xout252, xout253, xout254, xout255, xout256,
                yout1, yout2, yout3, yout4, yout5, yout6, yout7, yout8, yout9, yout10, yout11, yout12, yout13, yout14, yout15, yout16, yout17, yout18, yout19, yout20, yout21, yout22, yout23, yout24, yout25, yout26, yout27, yout28, yout29, yout30, yout31, yout32, yout33, yout34, yout35, yout36, yout37, yout38, yout39, yout40, yout41, yout42, yout43, yout44, yout45, yout46, yout47, yout48, yout49, yout50, yout51, yout52, yout53, yout54, yout55, yout56, yout57, yout58, yout59, yout60, yout61, yout62, yout63, yout64, yout65, yout66, yout67, yout68, yout69, yout70, yout71, yout72, yout73, yout74, yout75, yout76, yout77, yout78, yout79, yout80, yout81, yout82, yout83, yout84, yout85, yout86, yout87, yout88, yout89, yout90, yout91, yout92, yout93, yout94, yout95, yout96, yout97, yout98, yout99, yout100, yout101, yout102, yout103, yout104, yout105, yout106, yout107, yout108, yout109, yout110, yout111, yout112, yout113, yout114, yout115, yout116, yout117, yout118, yout119, yout120, yout121, yout122, yout123, yout124, yout125, yout126, yout127, yout128, yout129, yout130, yout131, yout132, yout133, yout134, yout135, yout136, yout137, yout138, yout139, yout140, yout141, yout142, yout143, yout144, yout145, yout146, yout147, yout148, yout149, yout150, yout151, yout152, yout153, yout154, yout155, yout156, yout157, yout158, yout159, yout160, yout161, yout162, yout163, yout164, yout165, yout166, yout167, yout168, yout169, yout170, yout171, yout172, yout173, yout174, yout175, yout176, yout177, yout178, yout179, yout180, yout181, yout182, yout183, yout184, yout185, yout186, yout187, yout188, yout189, yout190, yout191, yout192, yout193, yout194, yout195, yout196, yout197, yout198, yout199, yout200, yout201, yout202, yout203, yout204, yout205, yout206, yout207, yout208, yout209, yout210, yout211, yout212, yout213, yout214, yout215, yout216, yout217, yout218, yout219, yout220, yout221, yout222, yout223, yout224, yout225, yout226, yout227, yout228, yout229, yout230, yout231, yout232, yout233, yout234, yout235, yout236, yout237, yout238, yout239, yout240, yout241, yout242, yout243, yout244, yout245, yout246, yout247, yout248, yout249, yout250, yout251, yout252, yout253, yout254, yout255, yout256
        );




initial 
begin
    #100
    forever #5 clock = !clock;
end

initial
begin
   #100;
   
   		xin1=  1200;
		xin2 = 1200;
		xin3 = 1200;
		xin4 = 1200;
		xin5 = 1200;
		xin6 = 1200;
		xin7 = 1200;
		xin8 = 1200;
		xin9 = 1200;
		xin10 = 1200;
		xin11 = 1200;
	    xin12 = 1200;
	    xin13 = 1200;
	    xin14 = 1200;
	    xin15 = 1200;
	    xin16 = 1200;
	    xin17 = 3200;
end
endmodule
